/*
 * Copyright (c) 2003 Stephen Williams (steve@icarus.com)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 *
 *   $Id: process.v,v 1.1 2003/04/01 05:55:24 stevewilliams Exp $
 */

module process(output reg [7:0] upcounter,
	       output reg [7:0] downcounter,
	       input wire 	clk,
	       input wire 	reset);

   always @(posedge clk)
     if (reset)
       begin
	  upcounter <= 8'b0;
	  downcounter <= 8'b0;
       end
     else
       begin
	  upcounter <= upcounter + 1;
	  downcounter <= downcounter - 1;
       end

endmodule // process
